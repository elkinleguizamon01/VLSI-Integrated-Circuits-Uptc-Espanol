//AND gate in verilog

module ex2_and ( input logic a, b, 
            output logic y );
    assign y = a & b;
endmodule 
