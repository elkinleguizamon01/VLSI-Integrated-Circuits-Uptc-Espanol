//Or gate in verilog

module ex1 ( input logic a, b, 
            output logic y );
    assign y = a || b;
endmodule 
