//Or gate in verilog

module ex1_or ( input logic a, b, 
            output logic y );
    assign y = a || b;
endmodule 
